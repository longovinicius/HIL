--! \file		HIL_TOP.vhd
--!
--! \brief		
--!
--! \author		Vinícius de Carvalho Monteiro Longo (longo.vinicius@gmail.com)
--! \date       23-07-2025
--!
--! \version    1.0
--!
--! \copyright	Copyright (c) 2024 WEG - All Rights reserved.
--!
--! \note		Target devices : No specific target
--! \note		Tool versions  : No specific tool
--! \note		Dependencies   : No specific dependencies
--!
--! \ingroup	None
--! \warning	None
--!
--! \note		Revisions:
--!				- 1.0	23-07-2025	<longo.vinicius@gmail.com>
--!				First revision.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Solver_pkg.all;

entity HIL_TOP is
    port (
        SYSCLK_P                : in std_logic;
        SYSCLK_N                : in std_logic;
        PMOD6_PIN1_R            : in std_logic;
        
        GPIO_LED0               : out std_logic;
        GPIO_SW_C               : in std_logic;

        FT4232_B_UART_RX        : out std_logic;
        PMOD6_PIN3_R            : out std_logic
        --serial_data_out         : out std_logic_vector(0 to 4)
        
);
end entity HIL_TOP;

architecture arch of HIL_TOP is
    --------------------------------------------------------------------------
    -- Constants
    --------------------------------------------------------------------------
    constant CLK_FREQ           : integer := 200_000_000; 
    constant N_SS               : natural := 5;
    constant N_IN               : natural := 2;
    constant VDC_VOLTAGE        : integer := 400;
    constant RESET_TRSHD        : integer := 100;   
    constant START_PERIOD       : integer := 200; -- TODO: Investigar
    constant SERIAL_BAUD_RATE   : integer := 1_042_000;
    constant SERIAL_INTERVAL_US : integer := 200;
    
    constant L1                 : real := 1.0e-3;
    constant R1                 : real := 0.1;
    constant Cf                 : real := 3.3e-6;
    constant L2                 : real := 0.92e-3;
    constant R2                 : real := 0.1;
    constant Cd                 : real := 1.65e-6;
    constant Rd                 : real := 25.9;
    constant Ld                 : real := 5.1e-3;
    constant Ts                 : real := 1.0e-6;

    constant a00                : real := 1.0 - (R1/L1)*Ts; -- ok
    constant a03                : real := (-1.0/L1)*Ts; -- ok
    constant a13                : real := (1.0/Ld)*Ts;  -- ok
    constant a14                : real := (-1.0/Ld)*Ts; -- ok 
    constant a22                : real := 1.0 - (R2/L2)*Ts; -- ok
    constant a23                : real := (1.0/L2)*Ts; -- ok
    constant a30                : real := (1.0/Cf)*Ts; -- ok
    constant a31                : real := (-1.0/Cf)*Ts; -- ok
    constant a32                : real := (-1.0/Cf)*Ts; -- ok 
    constant a33                : real := 1.0 - (1.0/(Cf*Rd))*Ts; -- ok
    constant a34                : real := (1.0/(Cf*Rd))*Ts; -- ok
    constant a41                : real := (1.0/Cd)*Ts; -- ok
    constant a43                : real := (1.0/(Cd*Rd))*Ts; -- ok
    constant a44                : real := 1.0 - (1.0/(Cd*Rd))*Ts; -- ok
    constant b00                : real := (1.0/L1)*Ts;


    constant AMATRIX_C : matrix_fp_t(0 to N_SS - 1, 0 to N_SS - 1) := (
        (to_fp(a00), to_fp(0.0), to_fp(0.0), to_fp(a03), to_fp(0.0)),
        (to_fp(0.0), to_fp(1.0), to_fp(0.0), to_fp(a13), to_fp(a14)), 
        (to_fp(0.0), to_fp(0.0), to_fp(a22), to_fp(a23), to_fp(0.0)),
        (to_fp(a30), to_fp(a31), to_fp(a32), to_fp(a33), to_fp(a34)),
        (to_fp(0.0), to_fp(a41), to_fp(0.0), to_fp(a43), to_fp(a44))
    );

    constant BMATRIX_C : matrix_fp_t(0 to N_SS - 1, 0 to N_IN - 1) := (
        (to_fp(b00), to_fp(0.0)),
        (to_fp(0.0), to_fp(0.0)),
        (to_fp(0.0), to_fp(0.0)),
        (to_fp(0.0), to_fp(0.0)),
        (to_fp(0.0), to_fp(0.0))
    );

    constant XVEC_INITIAL_C : vector_fp_t(0 to N_SS - 1) := (
        to_fp(0.0), to_fp(0.0), to_fp(0.0), to_fp(0.0), to_fp(0.0)    
    );

    --------------------------------------------------------------------------
    -- Signals
    --------------------------------------------------------------------------
    signal sysclk_200mhz        : std_logic;
    signal reset_n              : std_logic := '0';
    signal reset_ctr            : unsigned(16 downto 0) := (others => '0');
    signal inverver_signal      : std_logic_vector(FP_TOTAL_BITS-1 downto 0);

    signal Xvec_current_o_sig   : vector_fp_t(0 to N_SS - 1);
    signal tx_out_sig           : std_logic_vector(0 to N_SS - 1);
    signal busy_o_sig           : std_logic;

    signal start_signal         : std_logic;
    signal start_ctr            : unsigned(26 downto 0) := (others => '0'); 
    signal Uvector              : vector_fp_t(0 to N_IN - 1) := (others => (others => '0') ); 

    signal pmod_sync_s1         : std_logic;
    signal pmod_sync_s2         : std_logic;

    signal serial_curr_L2_o     : std_logic; 

begin

    Synchronizer_Process: process (sysclk_200mhz)
    begin
        if rising_edge(sysclk_200mhz) then
            pmod_sync_s1 <= PMOD6_PIN1_R;
            pmod_sync_s2 <= pmod_sync_s1;
        end if;
    end process;

    --------------------------------------------------------------------------
    -- PLL
    --------------------------------------------------------------------------
    clock_gen_inst : entity work.clk_wiz_0
        port map(
            clk_in1_p => SYSCLK_P,
            clk_in1_n => SYSCLK_N,
            clk_out1  => sysclk_200mhz
        );

    --------------------------------------------------------------------------
    -- reset_n inicialization
    --------------------------------------------------------------------------
    process (sysclk_200mhz)
    begin
        if rising_edge(sysclk_200mhz) then
            if reset_ctr < RESET_TRSHD then
                reset_ctr <= reset_ctr + 1;
                reset_n   <= '0';
            else
                reset_n   <= '1';
            end if;
        end if;
    end process;

    --------------------------------------------------------------------------
    -- periodic start signal
    --------------------------------------------------------------------------
    process (sysclk_200mhz)
    begin
        if rising_edge(sysclk_200mhz) then
            if reset_n = '1' then
                if start_ctr < START_PERIOD - 1 then
                    start_ctr     <= start_ctr + 1;
                    start_signal  <= '0';
                else
                    start_ctr     <= (others => '0');
                    start_signal  <= '1'; 
                end if;
            else
                start_ctr     <= (others => '0');
                start_signal  <= '0';
            end if;
        end if;
    end process;

    --------------------------------------------------------------------------
    -- PWM to Voltage
    --------------------------------------------------------------------------
    PWMToVoltage_inst : entity work.PWMToVoltage
    generic map (
        VDC_VOLTAGE         => VDC_VOLTAGE,
        OUTPUT_BIT_WIDTH    => FP_TOTAL_BITS, 
        FP_FRACTION_BITS    => FP_FRACTION_BITS
    )
    port map (
        sysclk              => sysclk_200mhz,
        pwm_signal          => pmod_sync_s2,
        v_in                => inverver_signal
    );

    Uvector(0) <= inverver_signal;

    --------------------------------------------------------------------------
    -- LSM
    --------------------------------------------------------------------------
    LSM_inst : entity work.LinearSolver_Manager
    generic map (
        N_SS            => N_SS,
        N_IN            => N_IN
    )
    port map (
        sysclk         => sysclk_200mhz,
        reset_n        => reset_n,
        init_calc_i    => start_signal, 
        Amatrix_i      => AMATRIX_C,
        Bmatrix_i      => BMATRIX_C,
        Xvec_initial   => XVEC_INITIAL_C,
        Uvector_i      => Uvector,
        Xvec_current_o => Xvec_current_o_sig,
        busy_o         => busy_o_sig
    );

    --------------------------------------------------------------------------
    -- Serial Manager
    --------------------------------------------------------------------------
    -- SerialManager_gen : for index in 0 to N_SS-1 generate
    --     UUT_SerialManager : entity work.SerialManager
    --         generic map (
    --             CLK_FREQ          => CLK_FREQ,
    --             SEND_INTERVAL_US  => SERIAL_INTERVAL_US,
    --             BAUD_RATE         => SERIAL_BAUD_RATE
    --         )
    --         port map (
    --             sysclk            => sysclk_200mhz,
    --             reset_n           => reset_n,
    --             data_in_i         => Xvec_current_o_sig(index),
    --             tx_o              => tx_out_sig(index)
    --         );

    --     serial_data_out(index) <= tx_out_sig(index);
    -- end generate;

    UUT_SerialManager : entity work.SerialManager
        generic map (
            CLK_FREQ          => CLK_FREQ,
            SEND_INTERVAL_US  => SERIAL_INTERVAL_US,
            BAUD_RATE         => SERIAL_BAUD_RATE
        )
        port map (
            sysclk            => sysclk_200mhz,
            reset_n           => reset_n,
            data_in_i         => Xvec_current_o_sig(3),
            tx_o              => serial_curr_L2_o
        );
    --------------------------------------------------------------------------
    -- Output signals
    --------------------------------------------------------------------------
    GPIO_LED0 <= busy_o_sig;
    FT4232_B_UART_RX <= serial_curr_L2_o;
    PMOD6_PIN3_R <= serial_curr_L2_o;
    --------------------------------------------------------------------------
    -- ILA scope
    --------------------------------------------------------------------------
    -- chiscope_inst : entity work.ila_0
    --     port map(
    --         clk         => sysclk_200mhz,
    --         probe0      => start_signal,
    --         probe1      => pmod_sync_s2,               
    --         probe2      => busy_o_sig,                 
    --         probe3      => serial_curr_L2_o
    --     );

end architecture arch;